library verilog;
use verilog.vl_types.all;
entity contrl_vlg_vec_tst is
end contrl_vlg_vec_tst;
